//TODO
module tanh #(parameter ELEMENT_BITS = 8) (
		input logic		[ELEMENT_BITS-1:0]	data_in,
		output logic	[ELEMENT_BITS-1:0]	data_out
);
always_comb begin
	case(data_in)
		8'b00000000: data_out = 8'b00000000; // In = +0, 		Out = 0
		8'b00000001: data_out = 8'b00000001; // In = +0.015625, Out = 0.015625
		8'b00000010: data_out = 8'b00000010; // In = +0.03125,	Out = 0.03125
		8'b00000011: data_out = 8'b00000011; // In = +0.046875, Out = 0.046875
		8'b00000100: data_out = 8'b00000100; // In = +0.0625,	Out = 0.0625
		8'b00000101: data_out = 8'b00000101; // In = +0.078125,	Out = 0.078125
		8'b00000110: data_out = 8'b00000110; // In = +0.09375,	Out = 0.09375
		8'b00000111: data_out = 8'b00000111; // In = +0.109375,	Out = 0.109375
		8'b00001000: data_out = 8'b00001000; // In = +0.125,	Out = 0.125
		8'b00001001: data_out = 8'b00001001; // In = +0.140625,	Out = 0.140625
		8'b00001010: data_out = 8'b00001010; // In = +0.15625,	Out = 0.15625
		8'b00001011: data_out = 8'b00001011; // In = +0.171875,	Out = 0.171875
		8'b00001100: data_out = 8'b00001100; // In = +0.1875,	Out = 0.1875
		8'b00001101: data_out = 8'b00001101; // In = +0.203125,	Out = 0.203125
		8'b00001110: data_out = 8'b00001110; // In = +0.21875,	Out = 0.21875
		8'b00001111: data_out = 8'b00001111; // In = +0.234375,	Out = 0.234375
		8'b00010000: data_out = 8'b00010000; // In = +0.25,		Out = 0.25
		8'b00010001: data_out = 8'b00010001; // In = +0.265625,	Out = 0.265625
		8'b00010010: data_out = 8'b00010010; // In = +0.28125,	Out = 0.28125
		8'b00010011: data_out = 8'b00010011; // In = +0.296875,	Out = 0.296875
		8'b00010100: data_out = 8'b00010011; // In = +0.3125,	Out = 0.296875
		8'b00010101: data_out = 8'b00010100; // In = +0.328125,	Out = 0.3125
		8'b00010110: data_out = 8'b00010101; // In = +0.34375,	Out = 0.328125
		8'b00010111: data_out = 8'b00010110; // In = +0.359375,	Out = 0.34375
		8'b00011000: data_out = 8'b00010111; // In = +0.375,	Out = 0.359375
		8'b00011001: data_out = 8'b00011000; // In = +0.390625,	Out = 0.375
		8'b00011010: data_out = 8'b00011001; // In = +0.40625,	Out = 0.390625
		8'b00011011: data_out = 8'b00011010; // In = +0.421875,	Out = 0.40625
		8'b00011100: data_out = 8'b00011010; // In = +0.4375,	Out = 0.40625
		8'b00011101: data_out = 8'b00011011; // In = +0.453125,	Out = 0.421875
		8'b00011110: data_out = 8'b00011100; // In = +0.46875,	Out = 0.4375
		8'b00011111: data_out = 8'b00011101; // In = +0.484375,	Out = 0.453125
		8'b00100000: data_out = 8'b00011110; // In = +0.5,		Out = 0.46875
		8'b00100001: data_out = 8'b00011111; // In = +0.53125,	Out = 0.484375
		8'b00100010: data_out = 8'b00100000; // In = +0.5625,	Out = 0.5
		8'b00100011: data_out = 8'b00100001; // In = +0.59375,	Out = 0.53125
		8'b00100100: data_out = 8'b00100010; // In = +0.625,	Out = 0.5625
		8'b00100101: data_out = 8'b00100010; // In = +0.65625,	Out = 0.5625
		8'b00100110: data_out = 8'b00100011; // In = +0.6875,	Out = 0.59375
		8'b00100111: data_out = 8'b00100100; // In = +0.71875,	Out = 0.625
		8'b00101000: data_out = 8'b00100100; // In = +0.75,		Out = 0.625
		8'b00101001: data_out = 8'b00100101; // In = +0.78125,	Out = 0.65625
		8'b00101010: data_out = 8'b00100110; // In = +0.8125,	Out = 0.6875
		8'b00101011: data_out = 8'b00100110; // In = +0.84375,	Out = 0.6875
		8'b00101100: data_out = 8'b00100111; // In = +0.875,	Out = 0.71875
		8'b00101101: data_out = 8'b00100111; // In = +0.90625,	Out = 0.71875
		8'b00101110: data_out = 8'b00101000; // In = +0.9375,	Out = 0.75
		8'b00101111: data_out = 8'b00101000; // In = +0.96875,	Out = 0.75
		8'b00110000: data_out = 8'b00101000; // In = +1,		Out = 0.75
		8'b00110001: data_out = 8'b00101001; // In = +1.0625,	Out = 0.78125
		8'b00110010: data_out = 8'b00101010; // In = +1.125,	Out = 0.8125
		8'b00110011: data_out = 8'b00101010; // In = +1.1875,	Out = 0.8125
		8'b00110100: data_out = 8'b00101011; // In = +1.25,		Out = 0.84375
		8'b00110101: data_out = 8'b00101100; // In = +1.3125,	Out = 0.875
		8'b00110110: data_out = 8'b00101100; // In = +1.375,	Out = 0.875
		8'b00110111: data_out = 8'b00101101; // In = +1.4375,	Out = 0.90625
		8'b00111000: data_out = 8'b00101101; // In = +1.5,		Out = 0.90625
		8'b00111001: data_out = 8'b00101101; // In = +1.5625,	Out = 0.90625
		8'b00111010: data_out = 8'b00101110; // In = +1.625,	Out = 0.9375
		8'b00111011: data_out = 8'b00101110; // In = +1.6875,	Out = 0.9375
		8'b00111100: data_out = 8'b00101110; // In = +1.75,		Out = 0.9375
		8'b00111101: data_out = 8'b00101110; // In = +1.8125,	Out = 0.9375
		8'b00111110: data_out = 8'b00101111; // In = +1.875,	Out = 0.96875
		8'b00111111: data_out = 8'b00101111; // In = +1.9375,	Out = 0.96875
		8'b01000000: data_out = 8'b00101111; // In = +2,		Out = 0.96875
		8'b01000001: data_out = 8'b00101111; // In = +2.125, 	Out = 0.96875
		8'b01000010: data_out = 8'b00101111; // In = +2.25,	 	Out = 0.96875
		8'b01000011: data_out = 8'b00101111; // In = +2.375, 	Out = 0.96875
		8'b01000100: data_out = 8'b00110000; // In = +2.5, 	 	Out = 1 (clipped Here)
		8'b01000101: data_out = 8'b00110000; // In = +2.625, 	Out = 1
		8'b01000110: data_out = 8'b00110000; // In = +2.75,  	Out = 1
		8'b01000111: data_out = 8'b00110000; // In = +2.875, 	Out = 1
		8'b01001000: data_out = 8'b00110000; // In = +3.0,		Out = 1
		8'b01001001: data_out = 8'b00110000; // In = +3.125,	Out = 1
		8'b01001010: data_out = 8'b00110000; // In = +3.25,		Out = 1
		8'b01001011: data_out = 8'b00110000; // In = +3.375,	Out = 1
		8'b01001100: data_out = 8'b00110000; // In = +3.5,		Out = 1
		8'b01001101: data_out = 8'b00110000; // In = +3.625,	Out = 1
		8'b01001110: data_out = 8'b00110000; // In = +3.75,		Out = 1
		8'b01001111: data_out = 8'b00110000; // In = +3.875,	Out = 1
		8'b01010000: data_out = 8'b00110000; // In = +4.0,		Out = 1
		8'b01010001: data_out = 8'b00110000; // >4
		8'b01010010: data_out = 8'b00110000; // >4
		8'b01010011: data_out = 8'b00110000; // >4
		8'b01010100: data_out = 8'b00110000; // >4
		8'b01010101: data_out = 8'b00110000; // >4
		8'b01010110: data_out = 8'b00110000; // >4
		8'b01010111: data_out = 8'b00110000; // >4
		8'b01011000: data_out = 8'b00110000; // >4
		8'b01011001: data_out = 8'b00110000; // >4
		8'b01011010: data_out = 8'b00110000; // >4
		8'b01011011: data_out = 8'b00110000; // >4
		8'b01011100: data_out = 8'b00110000; // >4
		8'b01011101: data_out = 8'b00110000; // >4
		8'b01011110: data_out = 8'b00110000; // >4
		8'b01011111: data_out = 8'b00110000; // >4
		8'b01100000: data_out = 8'b00110000; // >4
		8'b01100001: data_out = 8'b00110000; // >4
		8'b01100010: data_out = 8'b00110000; // >4
		8'b01100011: data_out = 8'b00110000; // >4
		8'b01100100: data_out = 8'b00110000; // >4
		8'b01100101: data_out = 8'b00110000; // >4
		8'b01100110: data_out = 8'b00110000; // >4
		8'b01100111: data_out = 8'b00110000; // >4
		8'b01101000: data_out = 8'b00110000; // >4
		8'b01101001: data_out = 8'b00110000; // >4
		8'b01101010: data_out = 8'b00110000; // >4
		8'b01101011: data_out = 8'b00110000; // >4
		8'b01101100: data_out = 8'b00110000; // >4
		8'b01101101: data_out = 8'b00110000; // >4
		8'b01101110: data_out = 8'b00110000; // >4
		8'b01101111: data_out = 8'b00110000; // >4
		8'b01110000: data_out = 8'b00110000; // >4
		8'b01110001: data_out = 8'b00110000; // >4
		8'b01110010: data_out = 8'b00110000; // >4
		8'b01110011: data_out = 8'b00110000; // >4
		8'b01110100: data_out = 8'b00110000; // >4
		8'b01110101: data_out = 8'b00110000; // >4
		8'b01110110: data_out = 8'b00110000; // >4
		8'b01110111: data_out = 8'b00110000; // >4
		8'b01111000: data_out = 8'b00110000; // >4
		8'b01111001: data_out = 8'b00110000; // >4
		8'b01111010: data_out = 8'b00110000; // >4
		8'b01111011: data_out = 8'b00110000; // >4
		8'b01111100: data_out = 8'b00110000; // >4
		8'b01111101: data_out = 8'b00110000; // >4
		8'b01111110: data_out = 8'b00110000; // >4
		8'b01111111: data_out = 8'b00110000; // >4
		
		
		
		8'b10000000: data_out = 8'b10000000; // In = -0,		Out = 0
		8'b10000001: data_out = 8'b10000001; // In = -0.015625,	Out = -0.015625
		8'b10000010: data_out = 8'b10000010; // In = -0.03125,	Out = -0.03125
		8'b10000011: data_out = 8'b10000011; // In = -0.046875,	Out = -0.046875
		8'b10000100: data_out = 8'b10000100; // In = -0.0625,	Out = -0.0625
		8'b10000101: data_out = 8'b10000101; // In = -0.078125,	Out = -0.078125
		8'b10000110: data_out = 8'b10000110; // In = -0.09375,	Out = -0.09375
		8'b10000111: data_out = 8'b10000111; // In = -0.109375,	Out = -0.109375
		8'b10001000: data_out = 8'b10001000; // In = -0.125,	Out = -0.125
		8'b10001001: data_out = 8'b10001001; // In = -0.140625,	Out = -0.140625
		8'b10001010: data_out = 8'b10001010; // In = -0.15625,	Out = -0.15625
		8'b10001011: data_out = 8'b10001011; // In = -0.171875,	Out = -0.171875
		8'b10001100: data_out = 8'b10001100; // In = -0.1875,	Out = -0.1875
		8'b10001101: data_out = 8'b10001101; // In = -0.203125,	Out = -0.203125
		8'b10001110: data_out = 8'b10001110; // In = -0.21875,	Out = -0.21875
		8'b10001111: data_out = 8'b10001111; // In = -0.234375,	Out = -0.234375
		8'b10010000: data_out = 8'b10010000; // In = -0.25,		Out = -0.25
		8'b10010001: data_out = 8'b10010001; // In = -0.265625,	Out = -0.265625
		8'b10010010: data_out = 8'b10010010; // In = -0.28125,	Out = -0.28125
		8'b10010011: data_out = 8'b10010011; // In = -0.296875,	Out = -0.296875
		8'b10010100: data_out = 8'b10010011; // In = -0.3125,	Out = -0.296875
		8'b10010101: data_out = 8'b10010100; // In = -0.328125,	Out = -0.3125
		8'b10010110: data_out = 8'b10010101; // In = -0.34375,	Out = -0.328125
		8'b10010111: data_out = 8'b10010110; // In = -0.359375,	Out = -0.34375
		8'b10011000: data_out = 8'b10010111; // In = -0.375,	Out = -0.359375
		8'b10011001: data_out = 8'b10011000; // In = -0.390625,	Out = -0.375
		8'b10011010: data_out = 8'b10011001; // In = -0.40625,	Out = -0.390625
		8'b10011011: data_out = 8'b10011010; // In = -0.421875,	Out = -0.40625
		8'b10011100: data_out = 8'b10011010; // In = -0.4375,	Out = -0.40625
		8'b10011101: data_out = 8'b10011011; // In = -0.453125,	Out = -0.421875
		8'b10011110: data_out = 8'b10011100; // In = -0.46875,	Out = -0.4375
		8'b10011111: data_out = 8'b10011101; // In = -0.484375,	Out = -0.453125
		8'b10100000: data_out = 8'b10011110; // In = -0.5,		Out = -0.46875
		8'b10100001: data_out = 8'b10011111; // In = -0.53125,	Out = -0.484375
		8'b10100010: data_out = 8'b10100000; // In = -0.5625,	Out = -0.5
		8'b10100011: data_out = 8'b10100001; // In = -0.59375,	Out = -0.53125
		8'b10100100: data_out = 8'b10100010; // In = -0.625,	Out = -0.5625
		8'b10100101: data_out = 8'b10100010; // In = -0.65625,	Out = -0.5625
		8'b10100110: data_out = 8'b10100011; // In = -0.6875,	Out = -0.59375
		8'b10100111: data_out = 8'b10100100; // In = -0.71875,	Out = -0.625
		8'b10101000: data_out = 8'b10100100; // In = -0.75,		Out = -0.625
		8'b10101001: data_out = 8'b10100101; // In = -0.78125,	Out = -0.65625
		8'b10101010: data_out = 8'b10100110; // In = -0.8125,	Out = -0.6875
		8'b10101011: data_out = 8'b10100110; // In = -0.84375,	Out = -0.6875
		8'b10101100: data_out = 8'b10100111; // In = -0.875,	Out = -0.71875
		8'b10101101: data_out = 8'b10100111; // In = -0.90625,	Out = -0.71875
		8'b10101110: data_out = 8'b10101000; // In = -0.9375,	Out = -0.75
		8'b10101111: data_out = 8'b10101000; // In = -0.96875,	Out = -0.75
		8'b10110000: data_out = 8'b10101000; // In = -1.0,		Out = -0.75
		8'b10110001: data_out = 8'b10101001; // In = -1.0625,	Out = -0.0.78125
		8'b10110010: data_out = 8'b10101010; // In = -1.125,	Out = -0.8125
		8'b10110011: data_out = 8'b10101010; // In = -1.1875,	Out = -0.8125
		8'b10110100: data_out = 8'b10101011; // In = -1.25,		Out = -0.84375
		8'b10110101: data_out = 8'b10101100; // In = -1.3125,	Out = -0.875
		8'b10110110: data_out = 8'b10101100; // In = -1.375,	Out = -0.875
		8'b10110111: data_out = 8'b10101101; // In = -1.4375,	Out = -0.90625
		8'b10111000: data_out = 8'b10101101; // In = -1.5,		Out = -0.90625
		8'b10111001: data_out = 8'b10101101; // In = -1.5625,	Out = -0.90625
		8'b10111010: data_out = 8'b10101110; // In = -1.625,	Out = -0.9375
		8'b10111011: data_out = 8'b10101110; // In = -1.6875,	Out = -0.9375
		8'b10111100: data_out = 8'b10101110; // In = -1.75,		Out = -0.9375
		8'b10111101: data_out = 8'b10101110; // In = -1.8125,	Out = -0.9375
		8'b10111110: data_out = 8'b10101111; // In = -1.875,	Out = -0.96875
		8'b10111111: data_out = 8'b10101111; // In = -1.9375,	Out = -0.96875
		8'b11000000: data_out = 8'b10101111; // In = -2.0,		Out = -0.96875
		8'b11000001: data_out = 8'b10101111; // In = -2.125,	Out = -0.96875
		8'b11000010: data_out = 8'b10101111; // In = -2.25,		Out = -0.96875
		8'b11000011: data_out = 8'b10101111; // In = -2.375,	Out = -0.96875
		8'b11000100: data_out = 8'b10110000; // In = -2.5,		Out = -1 (clipped Here)
		8'b11000101: data_out = 8'b10110000; // In = -2.625,	Out = -1
		8'b11000110: data_out = 8'b10110000; // In = -2.75,		Out = -1
		8'b11000111: data_out = 8'b10110000; // In = -2.875,	Out = -1
		8'b11001000: data_out = 8'b10110000; // In = -3.0,		Out = -1
		8'b11001001: data_out = 8'b10110000; // In = -3.125,	Out = -1
		8'b11001010: data_out = 8'b10110000; // In = -3.25,		Out = -1
		8'b11001011: data_out = 8'b10110000; // In = -3.375,	Out = -1
		8'b11001100: data_out = 8'b10110000; // In = -3.5,		Out = -1
		8'b11001101: data_out = 8'b10110000; // In = -3.625,	Out = -1
		8'b11001110: data_out = 8'b10110000; // In = -3.75,		Out = -1
		8'b11001111: data_out = 8'b10110000; // In = -3.875,	Out = -1
		8'b11010000: data_out = 8'b10110000; // In = -4.0,		Out = -1
		8'b11010001: data_out = 8'b10110000; // <-4
		8'b11010010: data_out = 8'b10110000; // <-4
		8'b11010011: data_out = 8'b10110000; // <-4
		8'b11010100: data_out = 8'b10110000; // <-4
		8'b11010101: data_out = 8'b10110000; // <-4
		8'b11010110: data_out = 8'b10110000; // <-4
		8'b11010111: data_out = 8'b10110000; // <-4
		8'b11011000: data_out = 8'b10110000; // <-4
		8'b11011001: data_out = 8'b10110000; // <-4
		8'b11011010: data_out = 8'b10110000; // <-4
		8'b11011011: data_out = 8'b10110000; // <-4
		8'b11011100: data_out = 8'b10110000; // <-4
		8'b11011101: data_out = 8'b10110000; // <-4
		8'b11011110: data_out = 8'b10110000; // <-4
		8'b11011111: data_out = 8'b10110000; // <-4
		8'b11100000: data_out = 8'b10110000; // <-4
		8'b11100001: data_out = 8'b10110000; // <-4
		8'b11100010: data_out = 8'b10110000; // <-4
		8'b11100011: data_out = 8'b10110000; // <-4
		8'b11100100: data_out = 8'b10110000; // <-4
		8'b11100101: data_out = 8'b10110000; // <-4
		8'b11100110: data_out = 8'b10110000; // <-4
		8'b11100111: data_out = 8'b10110000; // <-4
		8'b11101000: data_out = 8'b10110000; // <-4
		8'b11101001: data_out = 8'b10110000; // <-4
		8'b11101010: data_out = 8'b10110000; // <-4
		8'b11101011: data_out = 8'b10110000; // <-4
		8'b11101100: data_out = 8'b10110000; // <-4
		8'b11101101: data_out = 8'b10110000; // <-4
		8'b11101110: data_out = 8'b10110000; // <-4
		8'b11101111: data_out = 8'b10110000; // <-4
		8'b11110000: data_out = 8'b10110000; // <-4
		8'b11110001: data_out = 8'b10110000; // <-4
		8'b11110010: data_out = 8'b10110000; // <-4
		8'b11110011: data_out = 8'b10110000; // <-4
		8'b11110100: data_out = 8'b10110000; // <-4
		8'b11110101: data_out = 8'b10110000; // <-4
		8'b11110110: data_out = 8'b10110000; // <-4
		8'b11110111: data_out = 8'b10110000; // <-4
		8'b11111000: data_out = 8'b10110000; // <-4
		8'b11111001: data_out = 8'b10110000; // <-4
		8'b11111010: data_out = 8'b10110000; // <-4
		8'b11111011: data_out = 8'b10110000; // <-4
		8'b11111100: data_out = 8'b10110000; // <-4
		8'b11111101: data_out = 8'b10110000; // <-4
		8'b11111110: data_out = 8'b10110000; // <-4
		8'b11111111: data_out = 8'b10110000; // <-4
        default: 	 data_out = 8'b10110000; // Default
	endcase
end
endmodule