
module mult_tb;

logic	[7:0]	in_a ;
logic	[7:0]	in_b ;
logic	[7:0]	res  ;

mult_top uut (.in_a(in_a),.in_b(in_b),.res(res)) ; 

initial begin
	in_a = 8'b00010101 ; //0.328125
	in_b = 8'b01000101 ; //2.625
	//res=(0.86132)10 ~= (0.875)10 = (0 010 1100)2
	#100
	in_a = 8'b00001000 ; //0.125
	in_b = 8'b01001001 ; //3.125
	//res=(0.390)10 ~= (0.390625)10 = (0 001 1001)2
	#100
	in_a = 8'b00101000 ; //0.75
	in_b = 8'b00101001 ; //0.78125
	//res=(0.585)10 ~= (0.59375)10 = (0 010 0011)2
	#100
	in_a = 8'b00111000 ; //1.5
	in_b = 8'b00101001 ; //0.78125
	//res=(1.171)10 ~= (1.1875)10 = (0 011 0011)2
	#100
	in_a = 8'b00101000 ; //0.75
	in_b = 8'b00111000 ; //1.5
	//res=(1.125)10 ~= (1.125)10 = (0 011 0010)2
	#100
	in_a = 8'b00001000 ; //0.125
	in_b = 8'b00010101 ; //0.328125
	//res=(0.0410)10 ~= (0.046875)10 = (0 000 0011)2
	#100
	in_a = 8'b00101000 ; //0.75
	in_b = 8'b00001000 ; //0.125
	//res=(0.09375)10 ~= (0.09375)10 = (0 000 0110)2
	#100
	in_a = 8'b00101000 ; //0.75
	in_b = 8'b01001001 ; //3.125
	//res=(2.34375)10 ~= (2.375)10 = (0 100 0011)2
	#100
	in_a = 8'b00010101 ; //0.328125
	in_b = 8'b00111000 ; //1.5
	//res=(0.4921875)10 ~= (0.5)10 = (0 010 0000)2
	#100
	in_a = 8'b00001000 ; //0.125
	in_b = 8'b00101001 ; //0.78125
	//res=(0.097656)10 ~= (0.09375)10 = (0 000 0110)2
	#100
	in_a = 8'b01101001 ; //3.125
	in_b = 8'b01101001 ; //3.125
	//res=(156.25)10 ~= (infty)10 = (0 111 0000)2
end

endmodule